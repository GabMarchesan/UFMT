library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity carry_adder is
  port( A, B: in STD_LOGIC_VECTOR(3 downto 0);
		   cin: in STD_LOGIC;
           S: out STD_LOGIC_VECTOR(3 downto 0);
		  cout: out STD_LOGIC
		  );
end carry_adder;

architecture synth of carry_adder is
    component fulladder is
        port(
            a, b, cin: in  STD_LOGIC;
            s, cout:   out STD_LOGIC
        );
    end component;

    signal cout1, cout2, cout3: STD_LOGIC;
begin

	FA1: fulladder port map( A(0), B(0), cin, S(0), cout1);
	FA2: fulladder port map( A(1), B(1), cout1, S(1), cout2);
	FA3: fulladder port map( A(2), B(2), cout2, S(2), cout3);
	FA4: fulladder port map( A(3), B(3), cout3, S(3), cout);
end synth;